--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

library work ;
use work.image_pack.all ;
use work.filter_pack.all ;
use work.blob_pack.all ;
use work.feature_pack.all ;
use work.graphic_pack.all ;
use work.interface_pack.all ;
use work.primitive_pack.all ;
use work.utils_pack.all ;

package hardcv_pack is


end hardcv_pack;

package body hardcv_pack is
 
end hardcv_pack;
